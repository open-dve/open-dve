`define odve_rand ( obj ) \
obj.user_randomize();