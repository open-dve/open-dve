module top;
    
    apb_if apb_if ();

    repeat (30) $display ("Hello world")
endmodule 
