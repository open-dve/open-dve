package odve_uart_agent_pkg;
    `include "odve_uart_item.sv"
    `include "odve_uart_driver.sv"
    `include "odve_uart_monitor.sv"
endpackage 