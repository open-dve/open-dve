module top;
    
    apb_if apb_if ();

    initial repeat (30) $display ("Hello world");
endmodule 
