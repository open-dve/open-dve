interface axi_if;
    
    
endinterface