interface odve_uart_if (
	input rx,
	output tx
	);
endinterface