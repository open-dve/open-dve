`ifndef __TEST_PKG_SV
`define __TEST_PKG_SV

package test_pkg;
    `include "uvm_macros.svh"
    import uvm_pkg::*;

    `include "read_test.sv"
endpackage  

`endif
