`ifndef ODVE_APB_SEQ_LIB_PKG__SV__
`define ODVE_APB_SEQ_LIB_PKG__SV__

package odve_apb_seq_lib_pkg ;
    `include "odve_apb_base_seq.sv"
    `include "odve_apb_read_seq.sv"
    `include "odve_apb_write_seq.sv"
endpackage 

`endif