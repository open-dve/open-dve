module dut (
    input clk, rst 
);
    
    initial repeat (1) $display ("Hi from DUT");
endmodule 
